typedef uvm_sequencer#(rd_tx) rd_sqr;