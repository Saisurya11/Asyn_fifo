typedef uvm_sequencer#(wr_tx) wr_sqr;